module ff_nnetwork(

)