module jn