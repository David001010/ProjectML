
module sys (
	clk_clk,
	reset_reset_n,
	uart_rxd,
	uart_txd);	

	input		clk_clk;
	input		reset_reset_n;
	input		uart_rxd;
	output		uart_txd;
endmodule
